d13 1
a13 1
// $Id: at_latch_h.v,v 1.1 2002/05/21 23:55:42 berndt Exp $
d27 1
a27 1
always @(negedge clk) begin
