
// $Id: j_rp01.v,v 1.1 2002/09/30 23:10:58 jeff Exp $

module j_rp01 (z);
   inout z;
   // supply0 vss;
   // nmos (z, z, vss);
   // trireg (medium) #(0.01, 0.01, 999999999) z;
endmodule
