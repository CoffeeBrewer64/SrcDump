a4 2
// XXX split into four module based on pinout;

d14 4
d74 8
d385 27
