
module rsp_lden32_f(ld_bar,clk,en_f);
input  [31:0] ld_bar;
input clk;
output [31:0] en_f;

or02d2 u00(.z(en_f[ 0]), .a1(ld_bar[ 0]), .a2(clk));
or02d2 u01(.z(en_f[ 1]), .a1(ld_bar[ 1]), .a2(clk));
or02d2 u02(.z(en_f[ 2]), .a1(ld_bar[ 2]), .a2(clk));
or02d2 u03(.z(en_f[ 3]), .a1(ld_bar[ 3]), .a2(clk));
or02d2 u04(.z(en_f[ 4]), .a1(ld_bar[ 4]), .a2(clk));
or02d2 u05(.z(en_f[ 5]), .a1(ld_bar[ 5]), .a2(clk));
or02d2 u06(.z(en_f[ 6]), .a1(ld_bar[ 6]), .a2(clk));
or02d2 u07(.z(en_f[ 7]), .a1(ld_bar[ 7]), .a2(clk));
or02d2 u08(.z(en_f[ 8]), .a1(ld_bar[ 8]), .a2(clk));
or02d2 u09(.z(en_f[ 9]), .a1(ld_bar[ 9]), .a2(clk));
or02d2 u10(.z(en_f[10]), .a1(ld_bar[10]), .a2(clk));
or02d2 u11(.z(en_f[11]), .a1(ld_bar[11]), .a2(clk));
or02d2 u12(.z(en_f[12]), .a1(ld_bar[12]), .a2(clk));
or02d2 u13(.z(en_f[13]), .a1(ld_bar[13]), .a2(clk));
or02d2 u14(.z(en_f[14]), .a1(ld_bar[14]), .a2(clk));
or02d2 u15(.z(en_f[15]), .a1(ld_bar[15]), .a2(clk));
or02d2 u16(.z(en_f[16]), .a1(ld_bar[16]), .a2(clk));
or02d2 u17(.z(en_f[17]), .a1(ld_bar[17]), .a2(clk));
or02d2 u18(.z(en_f[18]), .a1(ld_bar[18]), .a2(clk));
or02d2 u19(.z(en_f[19]), .a1(ld_bar[19]), .a2(clk));
or02d2 u20(.z(en_f[20]), .a1(ld_bar[20]), .a2(clk));
or02d2 u21(.z(en_f[21]), .a1(ld_bar[21]), .a2(clk));
or02d2 u22(.z(en_f[22]), .a1(ld_bar[22]), .a2(clk));
or02d2 u23(.z(en_f[23]), .a1(ld_bar[23]), .a2(clk));
or02d2 u24(.z(en_f[24]), .a1(ld_bar[24]), .a2(clk));
or02d2 u25(.z(en_f[25]), .a1(ld_bar[25]), .a2(clk));
or02d2 u26(.z(en_f[26]), .a1(ld_bar[26]), .a2(clk));
or02d2 u27(.z(en_f[27]), .a1(ld_bar[27]), .a2(clk));
or02d2 u28(.z(en_f[28]), .a1(ld_bar[28]), .a2(clk));
or02d2 u29(.z(en_f[29]), .a1(ld_bar[29]), .a2(clk));
or02d2 u30(.z(en_f[30]), .a1(ld_bar[30]), .a2(clk));
or02d2 u31(.z(en_f[31]), .a1(ld_bar[31]), .a2(clk));

endmodule
