d13 1
a13 1
// $Id: ram_bist_imem.v,v 1.1 2002/03/28 00:26:13 berndt Exp $
d166 1
a166 1
  always @(posedge clk or negedge reset_l)
d197 1
a197 1
  always @(posedge clk or negedge reset_l)
d233 1
a233 1
  always @(posedge clk or negedge reset_l)
