/**************************************************************************
 *                                                                        *
 *               Copyright (C) 1994, Silicon Graphics, Inc.               *
 *                                                                        *
 *  These coded instructions, statements, and computer programs  contain  *
 *  unpublished  proprietary  information of Silicon Graphics, Inc., and  *
 *  are protected by Federal copyright  law.  They  may not be disclosed  *
 *  to  third  parties  or copied or duplicated in any form, in whole or  *
 *  in part, without the prior written consent of Silicon Graphics, Inc.  *
 *                                                                        *
 *************************************************************************/
// $Id: inst_mux.v,v 1.1 2002/05/21 23:55:44 berndt Exp $

// inst_mux.v: 32-bit 8-input high-performance mux

`timescale 1ns / 10ps

module inst_mux (i0, i1, i2, i3, i4, i5, i6, i7, s0, s1, s2, z);

   input [31:0]		i0, i1, i2, i3, i4, i5, i6, i7;
   input 		s0, s1, s2;
   output [31:0]	z;


  mx81d1h mx81d1h_32_0 (.z(z[0]), .i0(i0[0]), .i1(i1[0]), .i2(i2[0]), .i3(i3[0]), .i4(i4[0]), .i5(i5[0]), .i6(i6[0]), .i7(i7[0]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_1 (.z(z[1]), .i0(i0[1]), .i1(i1[1]), .i2(i2[1]), .i3(i3[1]), .i4(i4[1]), .i5(i5[1]), .i6(i6[1]), .i7(i7[1]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_2 (.z(z[2]), .i0(i0[2]), .i1(i1[2]), .i2(i2[2]), .i3(i3[2]), .i4(i4[2]), .i5(i5[2]), .i6(i6[2]), .i7(i7[2]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_3 (.z(z[3]), .i0(i0[3]), .i1(i1[3]), .i2(i2[3]), .i3(i3[3]), .i4(i4[3]), .i5(i5[3]), .i6(i6[3]), .i7(i7[3]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_4 (.z(z[4]), .i0(i0[4]), .i1(i1[4]), .i2(i2[4]), .i3(i3[4]), .i4(i4[4]), .i5(i5[4]), .i6(i6[4]), .i7(i7[4]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_5 (.z(z[5]), .i0(i0[5]), .i1(i1[5]), .i2(i2[5]), .i3(i3[5]), .i4(i4[5]), .i5(i5[5]), .i6(i6[5]), .i7(i7[5]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_6 (.z(z[6]), .i0(i0[6]), .i1(i1[6]), .i2(i2[6]), .i3(i3[6]), .i4(i4[6]), .i5(i5[6]), .i6(i6[6]), .i7(i7[6]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_7 (.z(z[7]), .i0(i0[7]), .i1(i1[7]), .i2(i2[7]), .i3(i3[7]), .i4(i4[7]), .i5(i5[7]), .i6(i6[7]), .i7(i7[7]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_8 (.z(z[8]), .i0(i0[8]), .i1(i1[8]), .i2(i2[8]), .i3(i3[8]), .i4(i4[8]), .i5(i5[8]), .i6(i6[8]), .i7(i7[8]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_9 (.z(z[9]), .i0(i0[9]), .i1(i1[9]), .i2(i2[9]), .i3(i3[9]), .i4(i4[9]), .i5(i5[9]), .i6(i6[9]), .i7(i7[9]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_10 (.z(z[10]), .i0(i0[10]), .i1(i1[10]), .i2(i2[10]), .i3(i3[10]), .i4(i4[10]), .i5(i5[10]), .i6(i6[10]), .i7(i7[10]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_11 (.z(z[11]), .i0(i0[11]), .i1(i1[11]), .i2(i2[11]), .i3(i3[11]), .i4(i4[11]), .i5(i5[11]), .i6(i6[11]), .i7(i7[11]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_12 (.z(z[12]), .i0(i0[12]), .i1(i1[12]), .i2(i2[12]), .i3(i3[12]), .i4(i4[12]), .i5(i5[12]), .i6(i6[12]), .i7(i7[12]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_13 (.z(z[13]), .i0(i0[13]), .i1(i1[13]), .i2(i2[13]), .i3(i3[13]), .i4(i4[13]), .i5(i5[13]), .i6(i6[13]), .i7(i7[13]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_14 (.z(z[14]), .i0(i0[14]), .i1(i1[14]), .i2(i2[14]), .i3(i3[14]), .i4(i4[14]), .i5(i5[14]), .i6(i6[14]), .i7(i7[14]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_15 (.z(z[15]), .i0(i0[15]), .i1(i1[15]), .i2(i2[15]), .i3(i3[15]), .i4(i4[15]), .i5(i5[15]), .i6(i6[15]), .i7(i7[15]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_16 (.z(z[16]), .i0(i0[16]), .i1(i1[16]), .i2(i2[16]), .i3(i3[16]), .i4(i4[16]), .i5(i5[16]), .i6(i6[16]), .i7(i7[16]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_17 (.z(z[17]), .i0(i0[17]), .i1(i1[17]), .i2(i2[17]), .i3(i3[17]), .i4(i4[17]), .i5(i5[17]), .i6(i6[17]), .i7(i7[17]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_18 (.z(z[18]), .i0(i0[18]), .i1(i1[18]), .i2(i2[18]), .i3(i3[18]), .i4(i4[18]), .i5(i5[18]), .i6(i6[18]), .i7(i7[18]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_19 (.z(z[19]), .i0(i0[19]), .i1(i1[19]), .i2(i2[19]), .i3(i3[19]), .i4(i4[19]), .i5(i5[19]), .i6(i6[19]), .i7(i7[19]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_20 (.z(z[20]), .i0(i0[20]), .i1(i1[20]), .i2(i2[20]), .i3(i3[20]), .i4(i4[20]), .i5(i5[20]), .i6(i6[20]), .i7(i7[20]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_21 (.z(z[21]), .i0(i0[21]), .i1(i1[21]), .i2(i2[21]), .i3(i3[21]), .i4(i4[21]), .i5(i5[21]), .i6(i6[21]), .i7(i7[21]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_22 (.z(z[22]), .i0(i0[22]), .i1(i1[22]), .i2(i2[22]), .i3(i3[22]), .i4(i4[22]), .i5(i5[22]), .i6(i6[22]), .i7(i7[22]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_23 (.z(z[23]), .i0(i0[23]), .i1(i1[23]), .i2(i2[23]), .i3(i3[23]), .i4(i4[23]), .i5(i5[23]), .i6(i6[23]), .i7(i7[23]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_24 (.z(z[24]), .i0(i0[24]), .i1(i1[24]), .i2(i2[24]), .i3(i3[24]), .i4(i4[24]), .i5(i5[24]), .i6(i6[24]), .i7(i7[24]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_25 (.z(z[25]), .i0(i0[25]), .i1(i1[25]), .i2(i2[25]), .i3(i3[25]), .i4(i4[25]), .i5(i5[25]), .i6(i6[25]), .i7(i7[25]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_26 (.z(z[26]), .i0(i0[26]), .i1(i1[26]), .i2(i2[26]), .i3(i3[26]), .i4(i4[26]), .i5(i5[26]), .i6(i6[26]), .i7(i7[26]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_27 (.z(z[27]), .i0(i0[27]), .i1(i1[27]), .i2(i2[27]), .i3(i3[27]), .i4(i4[27]), .i5(i5[27]), .i6(i6[27]), .i7(i7[27]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_28 (.z(z[28]), .i0(i0[28]), .i1(i1[28]), .i2(i2[28]), .i3(i3[28]), .i4(i4[28]), .i5(i5[28]), .i6(i6[28]), .i7(i7[28]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_29 (.z(z[29]), .i0(i0[29]), .i1(i1[29]), .i2(i2[29]), .i3(i3[29]), .i4(i4[29]), .i5(i5[29]), .i6(i6[29]), .i7(i7[29]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_30 (.z(z[30]), .i0(i0[30]), .i1(i1[30]), .i2(i2[30]), .i3(i3[30]), .i4(i4[30]), .i5(i5[30]), .i6(i6[30]), .i7(i7[30]), .s0(s0), .s1(s1), .s2(s2)); 
  mx81d1h mx81d1h_32_31 (.z(z[31]), .i0(i0[31]), .i1(i1[31]), .i2(i2[31]), .i3(i3[31]), .i4(i4[31]), .i5(i5[31]), .i6(i6[31]), .i7(i7[31]), .s0(s0), .s1(s1), .s2(s2)); 

endmodule
