
// generally useful parameters
parameter
   LOW				= 1'b0,
   HIGH				= 1'b1;
  //  FLOAT			= 1'bz,
  //  UNKNOWN			= 1'bx;

// SysAD bus widths
// parameter SYS_AD_SIZE		= 32;
// parameter SYS_CMD_SIZE		= 5;
// parameter SYS_CMD_BLOCK_SIZE	= 2;

// SysCMD command bit definitions
// parameter
	// SYS_CMD_DATA		= 4,
	// SYS_CMD_WRITE		= 3,
	// SYS_CMD_BLOCK		= 2,
	// SYS_CMD_SIZE_START 	= 1,
	// SYS_CMD_SIZE_END	= 0,
	// SYS_CMD_MORE 		= 3,
	// SYS_CMD_ERROR		= 1;

// SysCMD word definitions
// parameter SYS_CMD_WRITE_WORD	= 5'b01000;
// parameter SYS_CMD_READ_WORD	= 5'b00000;
// parameter SYS_CMD_WRITE_BLOCK	= 5'b01100;
// parameter SYS_CMD_READ_BLOCK	= 5'b00100;
// parameter SYS_CMD_DATA_NEXT	= 5'b11000;
// parameter SYS_CMD_DATA_LAST	= 5'b10000;

// AD16 bus widths
// parameter AD16_DATA_SIZE	= 16;

// vbus bus widths
// parameter VBUS_DATA_SIZE	= 7;

// Rambus definitions
// parameter RAMBUS_DATA_SIZE	= 9;
