d13 1
a13 1
// $Id: ms_debug.v,v 1.1 2002/05/21 23:55:43 berndt Exp $
d123 1
a123 1
always @(posedge clock or negedge reset_l) begin
