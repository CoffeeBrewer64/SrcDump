d2 1
a2 1
// $Id: j_dfctnb.v,v 1.4 2002/11/13 01:38:38 rws Exp $
d12 1
a12 1
   always @ (posedge cp or negedge cdn) begin
