module div_rom(clk, oe, a, out);

input clk, oe;
input [9:0] a;
output [15:0] out;

endmodule
