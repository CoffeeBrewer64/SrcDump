d13 1
a13 1
// $Id: ram_bist_tmem.v,v 1.1 2002/03/28 00:26:14 berndt Exp $
d248 1
a248 1
  always @(posedge clk or negedge reset_l)
d279 1
a279 1
  always @(posedge clk or negedge reset_l)
d314 1
a314 1
  always @(posedge clk or negedge reset_l)
