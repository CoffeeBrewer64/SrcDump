d27 1
a27 1
always @(posedge clk) begin
