module tmem_driver(tmem_data_out, tmem_enable, tmem_data);

input [63:0] tmem_data_out;
input tmem_enable;
output [63:0] tmem_data;

assign tmem_data = tmem_enable ? tmem_data_out : {64{1'bz}};

// nt01d3 b0 (.i(tmem_data_out[0]), .z(tmem_data[0]), .oe(tmem_enable));
// nt01d3 b1 (.i(tmem_data_out[1]), .z(tmem_data[1]), .oe(tmem_enable));
// nt01d3 b2 (.i(tmem_data_out[2]), .z(tmem_data[2]), .oe(tmem_enable));
// nt01d3 b3 (.i(tmem_data_out[3]), .z(tmem_data[3]), .oe(tmem_enable));
// nt01d3 b4 (.i(tmem_data_out[4]), .z(tmem_data[4]), .oe(tmem_enable));
// nt01d3 b5 (.i(tmem_data_out[5]), .z(tmem_data[5]), .oe(tmem_enable));
// nt01d3 b6 (.i(tmem_data_out[6]), .z(tmem_data[6]), .oe(tmem_enable));
// nt01d3 b7 (.i(tmem_data_out[7]), .z(tmem_data[7]), .oe(tmem_enable));
// nt01d3 b8 (.i(tmem_data_out[8]), .z(tmem_data[8]), .oe(tmem_enable));
// nt01d3 b9 (.i(tmem_data_out[9]), .z(tmem_data[9]), .oe(tmem_enable));
// nt01d3 b10 (.i(tmem_data_out[10]), .z(tmem_data[10]), .oe(tmem_enable));
// nt01d3 b11 (.i(tmem_data_out[11]), .z(tmem_data[11]), .oe(tmem_enable));
// nt01d3 b12 (.i(tmem_data_out[12]), .z(tmem_data[12]), .oe(tmem_enable));
// nt01d3 b13 (.i(tmem_data_out[13]), .z(tmem_data[13]), .oe(tmem_enable));
// nt01d3 b14 (.i(tmem_data_out[14]), .z(tmem_data[14]), .oe(tmem_enable));
// nt01d3 b15 (.i(tmem_data_out[15]), .z(tmem_data[15]), .oe(tmem_enable));
// nt01d3 b16 (.i(tmem_data_out[16]), .z(tmem_data[16]), .oe(tmem_enable));
// nt01d3 b17 (.i(tmem_data_out[17]), .z(tmem_data[17]), .oe(tmem_enable));
// nt01d3 b18 (.i(tmem_data_out[18]), .z(tmem_data[18]), .oe(tmem_enable));
// nt01d3 b19 (.i(tmem_data_out[19]), .z(tmem_data[19]), .oe(tmem_enable));
// nt01d3 b20 (.i(tmem_data_out[20]), .z(tmem_data[20]), .oe(tmem_enable));
// nt01d3 b21 (.i(tmem_data_out[21]), .z(tmem_data[21]), .oe(tmem_enable));
// nt01d3 b22 (.i(tmem_data_out[22]), .z(tmem_data[22]), .oe(tmem_enable));
// nt01d3 b23 (.i(tmem_data_out[23]), .z(tmem_data[23]), .oe(tmem_enable));
// nt01d3 b24 (.i(tmem_data_out[24]), .z(tmem_data[24]), .oe(tmem_enable));
// nt01d3 b25 (.i(tmem_data_out[25]), .z(tmem_data[25]), .oe(tmem_enable));
// nt01d3 b26 (.i(tmem_data_out[26]), .z(tmem_data[26]), .oe(tmem_enable));
// nt01d3 b27 (.i(tmem_data_out[27]), .z(tmem_data[27]), .oe(tmem_enable));
// nt01d3 b28 (.i(tmem_data_out[28]), .z(tmem_data[28]), .oe(tmem_enable));
// nt01d3 b29 (.i(tmem_data_out[29]), .z(tmem_data[29]), .oe(tmem_enable));
// nt01d3 b30 (.i(tmem_data_out[30]), .z(tmem_data[30]), .oe(tmem_enable));
// nt01d3 b31 (.i(tmem_data_out[31]), .z(tmem_data[31]), .oe(tmem_enable));
// nt01d3 b32 (.i(tmem_data_out[32]), .z(tmem_data[32]), .oe(tmem_enable));
// nt01d3 b33 (.i(tmem_data_out[33]), .z(tmem_data[33]), .oe(tmem_enable));
// nt01d3 b34 (.i(tmem_data_out[34]), .z(tmem_data[34]), .oe(tmem_enable));
// nt01d3 b35 (.i(tmem_data_out[35]), .z(tmem_data[35]), .oe(tmem_enable));
// nt01d3 b36 (.i(tmem_data_out[36]), .z(tmem_data[36]), .oe(tmem_enable));
// nt01d3 b37 (.i(tmem_data_out[37]), .z(tmem_data[37]), .oe(tmem_enable));
// nt01d3 b38 (.i(tmem_data_out[38]), .z(tmem_data[38]), .oe(tmem_enable));
// nt01d3 b39 (.i(tmem_data_out[39]), .z(tmem_data[39]), .oe(tmem_enable));
// nt01d3 b40 (.i(tmem_data_out[40]), .z(tmem_data[40]), .oe(tmem_enable));
// nt01d3 b41 (.i(tmem_data_out[41]), .z(tmem_data[41]), .oe(tmem_enable));
// nt01d3 b42 (.i(tmem_data_out[42]), .z(tmem_data[42]), .oe(tmem_enable));
// nt01d3 b43 (.i(tmem_data_out[43]), .z(tmem_data[43]), .oe(tmem_enable));
// nt01d3 b44 (.i(tmem_data_out[44]), .z(tmem_data[44]), .oe(tmem_enable));
// nt01d3 b45 (.i(tmem_data_out[45]), .z(tmem_data[45]), .oe(tmem_enable));
// nt01d3 b46 (.i(tmem_data_out[46]), .z(tmem_data[46]), .oe(tmem_enable));
// nt01d3 b47 (.i(tmem_data_out[47]), .z(tmem_data[47]), .oe(tmem_enable));
// nt01d3 b48 (.i(tmem_data_out[48]), .z(tmem_data[48]), .oe(tmem_enable));
// nt01d3 b49 (.i(tmem_data_out[49]), .z(tmem_data[49]), .oe(tmem_enable));
// nt01d3 b50 (.i(tmem_data_out[50]), .z(tmem_data[50]), .oe(tmem_enable));
// nt01d3 b51 (.i(tmem_data_out[51]), .z(tmem_data[51]), .oe(tmem_enable));
// nt01d3 b52 (.i(tmem_data_out[52]), .z(tmem_data[52]), .oe(tmem_enable));
// nt01d3 b53 (.i(tmem_data_out[53]), .z(tmem_data[53]), .oe(tmem_enable));
// nt01d3 b54 (.i(tmem_data_out[54]), .z(tmem_data[54]), .oe(tmem_enable));
// nt01d3 b55 (.i(tmem_data_out[55]), .z(tmem_data[55]), .oe(tmem_enable));
// nt01d3 b56 (.i(tmem_data_out[56]), .z(tmem_data[56]), .oe(tmem_enable));
// nt01d3 b57 (.i(tmem_data_out[57]), .z(tmem_data[57]), .oe(tmem_enable));
// nt01d3 b58 (.i(tmem_data_out[58]), .z(tmem_data[58]), .oe(tmem_enable));
// nt01d3 b59 (.i(tmem_data_out[59]), .z(tmem_data[59]), .oe(tmem_enable));
// nt01d3 b60 (.i(tmem_data_out[60]), .z(tmem_data[60]), .oe(tmem_enable));
// nt01d3 b61 (.i(tmem_data_out[61]), .z(tmem_data[61]), .oe(tmem_enable));
// nt01d3 b62 (.i(tmem_data_out[62]), .z(tmem_data[62]), .oe(tmem_enable));
// nt01d3 b63 (.i(tmem_data_out[63]), .z(tmem_data[63]), .oe(tmem_enable));

endmodule
