d2 1
a2 1
// $Id: j_dfptnb.v,v 1.3 2002/11/13 01:38:38 rws Exp $
d12 1
a12 1
   always @ (posedge cp or negedge sdn) begin
